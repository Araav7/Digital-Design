`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// National University of Singapore
// Department of Electrical and Computer Engineering
// EE2026 Digital Design
// AY1819 Semester 1
// Project: Voice Scope
//////////////////////////////////////////////////////////////////////////////////

module Voice_Scope_TOP(
    input CLK,
    input [9:0]sw,
    input [4:0]btn,
    
    input  J_MIC3_Pin3,   // PmodMIC3 audio input data (serial)
    output J_MIC3_Pin1,   // PmodMIC3 chip select, 20kHz sampling clock
    output J_MIC3_Pin4,   // PmodMIC3 serial clock (generated by module VoiceCapturer.v)
   
    output [3:0] VGA_RED,    // RGB outputs to VGA connector (4 bits per channel gives 4096 possible colors)
    output [3:0] VGA_GREEN,
    output [3:0] VGA_BLUE,
    
    output VGA_VS,          // horizontal & vertical sync outputs to VGA connector
    output VGA_HS,
    output [11:0]led,
    output [3:0]an,
    output [6:0]seg
    
    );


      
       
//-----------------------------------------------------------------------------
//                  STUDENT A - MIC
//-----------------------------------------------------------------------------

       
                 
    wire clk1;
    wire [11:0]sample;
    wire [11:0]volume;
    wire [9:0]sample_max;
    
// Please create a clock divider module to generate a 20kHz clock signal. 
// Instantiate it below
    
    
    clk_div clock (CLK, clk1);
   
       
// Please instantiate the voice capturer module below
   


    Voice_Capturer capture (CLK, clk1, J_MIC3_Pin3, J_MIC3_Pin1, J_MIC3_Pin4, sample);
    indicator leds (CLK, sample, volume, sample_max);
    segments segs (CLK, volume, an, seg);
    assign led = volume;


//-----------------------------------------------------------------------------
//                  STUDENT B - VGA
//-----------------------------------------------------------------------------

    wire [9:0]ramp_sample;
    
    TestWave_Gen test (clk1, ramp_sample);

    wire [11:0] VGA_HORZ_COORD;
    wire [11:0] VGA_VERT_COORD; 
    wire [1:0] state;
    
// Please instantiate the background drawing module below   
    wire [3:0] VGA_Red_grid;
    wire [3:0] VGA_Green_grid;
    wire [3:0] VGA_Blue_grid;
   Draw_Background background (clk1, btn, sw, VGA_HORZ_COORD, VGA_VERT_COORD, VGA_Red_grid, VGA_Green_grid,
                            VGA_Blue_grid, state);
                            
// Please instantiate the waveform drawer module below
    
    wire [3:0] VGA_Red_waveform;
    wire [3:0] VGA_Green_waveform;
    wire [3:0] VGA_Blue_waveform;
    wire [9:0] wave_sample;
    
    assign wave_sample = (sw[4]) ? ramp_sample : sample[11:2];
    
    Draw_Waveform draw (state, btn[0], btn[1], btn[2], btn[3], sw, clk1, sample_max, wave_sample, VGA_HORZ_COORD, VGA_VERT_COORD, VGA_Red_waveform, VGA_Green_waveform,
                        VGA_Blue_waveform);
    

    
// Please instantiate the VGA display module below     
     
    VGA_DISPLAY display (CLK, VGA_Red_waveform, VGA_Green_waveform, VGA_Blue_waveform, VGA_Red_grid, VGA_Green_grid,
                         VGA_Blue_grid, VGA_HORZ_COORD, VGA_VERT_COORD, VGA_RED, VGA_GREEN, VGA_BLUE, VGA_VS, VGA_HS
    );
     
     
     
                    
endmodule
